
int no_of_pkts=100;
static int error=0;

